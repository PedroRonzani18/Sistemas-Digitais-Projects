/*
Nomes: Pedro Augusto, Tulio Horta
Projeto: somador geral
Data: 29/09/2022
*/

module somador (A,B,TE,S,TS);

	input A,B,TE;
	output S,TS;
	
endmodule