module decod(E,S);

	input [0:3]E;
	output [0:6]S;
	 
	//assign S[0] = (~E[0] & ~E[1] & ~E[2] &  E[3]) | (~E[0] & E[1] & ~E[2] & ~E[3]);
	//assign S[1] = (~E[0] &  E[1] & ~E[2] &  E[3]) | (~E[0] & E[1] &  E[2] & ~E[3]);
	//assign S[3] = (~E[0] & ~E[1] & ~E[2] &  E[3]) | (~E[0] & E[1] & ~E[2] & ~E[3]) | (~E[0] & E[1] & E[2] &  E[3]);
	//assign S[4] = E[3] | E[1] & E[2] & ~E[3] 
	
	
	assign S[0] = ( E[1] & ~E[2] &  ~E[3]) | (~E[0] & ~E[1] & ~E[2] & E[3]);
	assign S[1] = ( E[1] & ~E[2] &  E[3]) | ( E[1] &  E[2] & ~E[3]);
	assign S[2] = (~E[0] & ~E[1] &  E[2] & ~E[3]);
	assign S[3] = (~E[0] & ~E[1] & ~E[2] &  E[3]) | (E[1] & ~E[2] & ~E[3]) | (E[1] & E[2] &  E[3]);
	assign S[4] = ( E[3]) | (E[1] & ~E[2]);
	assign S[5] = ( E[2] & E[3]) | (~E[0] & ~E[1] & E[3]) | (~E[0] & ~E[1] & E[2]);
	assign S[6] = (~E[0] & ~E[1] & ~E[2]) | (E[1] & E[2] & E[3]);
	
endmodule